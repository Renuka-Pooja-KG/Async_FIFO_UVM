class base_test extends uvm_test;
  `uvm_component_utils(base_test)

  env m_env;
  write_base_sequence wseq;
  read_base_sequence rseq;

  function new(string name = "base_test", uvm_component parent = null);
    super.new(name, parent);
  endfunction

  function void build_phase(uvm_phase phase);
    super.build_phase(phase);
    m_env = env::type_id::create("m_env", this);
    wseq = write_base_sequence::type_id::create("wseq");
    rseq = read_base_sequence::type_id::create("rseq");
    `uvm_info(get_type_name(), "Base test build_phase completed", UVM_LOW)
  endfunction

  function void end_of_elaboration_phase(uvm_phase phase);
    super.end_of_elaboration_phase(phase);
    uvm_top.print_topology();
    `uvm_info(get_type_name(), "Base test end_of_elaboration_phase completed", UVM_LOW)
  endfunction

  task run_phase(uvm_phase phase);
    phase.raise_objection(this);
    
    // Configure scoreboard for data integrity priority mode
    configure_scoreboard_for_test();
    
    fork
      // Sequence starting should be done in derived tests
      wseq.start(m_env.m_write_agent.m_sequencer);
      rseq.start(m_env.m_read_agent.m_sequencer);
    join
    
    // Get and report data integrity statistics
    report_data_integrity_stats();
    
    `uvm_info(get_type_name(), "Base test run_phase - sequences should be applied in derived tests", UVM_LOW)
    phase.drop_objection(this);
  endtask
  
  // Function to configure scoreboard settings for different test types
  function void configure_scoreboard_for_test();
    // Default configuration: Enable data integrity priority and level mismatch tolerance
    m_env.m_scoreboard.set_data_integrity_priority(1'b1);
    m_env.m_scoreboard.set_level_mismatch_tolerance(1'b1);
    
    // Configure parameters based on test type
    configure_scoreboard_parameters();
    
    // Configure tolerance settings based on test type
    configure_scoreboard_tolerance();
    
    `uvm_info(get_type_name(), "Scoreboard configured for data integrity priority mode", UVM_MEDIUM)
  endfunction
  
  // Function to configure scoreboard parameters based on test type
  function void configure_scoreboard_parameters();
    // Default parameters
    int soft_reset_val = 3;  // Default SOFT_RESET value
    int sync_stage_val = 2;  // Default SYNC_STAGE value
    
    // Override parameters based on test type
    case (get_type_name())
      "sync_stage_3_test": begin
        sync_stage_val = 3;
        `uvm_info(get_type_name(), "Configuring scoreboard for SYNC_STAGE=3", UVM_MEDIUM)
      end
      "soft_reset_test": begin
        soft_reset_val = 3;
        `uvm_info(get_type_name(), "Configuring scoreboard for SOFT_RESET=3", UVM_MEDIUM)
      end
      "soft_reset_test_0": begin
        soft_reset_val = 0;
        `uvm_info(get_type_name(), "Configuring scoreboard for SOFT_RESET=0", UVM_MEDIUM)
      end
      "soft_reset_test_1": begin
        soft_reset_val = 1;
        `uvm_info(get_type_name(), "Configuring scoreboard for SOFT_RESET=1", UVM_MEDIUM)
      end
      "soft_reset_test_2": begin
        soft_reset_val = 2;
        `uvm_info(get_type_name(), "Configuring scoreboard for SOFT_RESET=2", UVM_MEDIUM)
      end
      default: begin
        // Use default values
        `uvm_info(get_type_name(), "Using default scoreboard parameters", UVM_MEDIUM)
      end
    endcase
    
    // Set the parameters in the scoreboard
    m_env.m_scoreboard.set_soft_reset_param(soft_reset_val);
    m_env.m_scoreboard.set_sync_stage_param(sync_stage_val);
    
    `uvm_info(get_type_name(), $sformatf("Scoreboard parameters configured: SOFT_RESET=%0d, SYNC_STAGE=%0d", soft_reset_val, sync_stage_val), UVM_MEDIUM)
  endfunction
  
  // Function to configure scoreboard tolerance settings based on test type
  function void configure_scoreboard_tolerance();
    // Default tolerance settings
    m_env.m_scoreboard.set_underflow_tolerance(1'b1);
    m_env.m_scoreboard.set_write_count_tolerance(1'b1);
    
    // Configure tolerance based on test type
    case (get_type_name())
      "sync_stage_3_test": begin
        // Enable write count tolerance for SYNC_STAGE=3 due to increased sync delays
        m_env.m_scoreboard.set_write_count_tolerance(1'b1);
        `uvm_info(get_type_name(), "Write count tolerance enabled for SYNC_STAGE=3", UVM_MEDIUM)
      end
      "soft_reset_test", "soft_reset_test_0", "soft_reset_test_1", "soft_reset_test_2": begin
        // Enable tolerance for soft reset tests
        m_env.m_scoreboard.set_write_count_tolerance(1'b1);
        m_env.m_scoreboard.set_reset_scenario_mode(1'b1);
        `uvm_info(get_type_name(), "Tolerance enabled for soft reset test", UVM_MEDIUM)
      end
      default: begin
        // Use default tolerance settings
        `uvm_info(get_type_name(), "Using default tolerance settings", UVM_MEDIUM)
      end
    endcase
  endfunction
  
  // Function to get and report data integrity statistics
  function void report_data_integrity_stats();
    int total_ops, sim_ops, errors;
    m_env.m_scoreboard.get_data_integrity_stats(total_ops, sim_ops, errors);
    `uvm_info(get_type_name(), $sformatf("Data Integrity Statistics: Total_Ops=%0d, Simultaneous_Ops=%0d, Errors=%0d", total_ops, sim_ops, errors), UVM_LOW)
  endfunction
endclass 