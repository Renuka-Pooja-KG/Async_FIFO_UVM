class scoreboard extends uvm_scoreboard;
    `uvm_component_utils(scoreboard)

    uvm_analysis_export #(write_sequence_item) write_export;
    uvm_analysis_export #(read_sequence_item)  read_export;

    uvm_tlm_analysis_fifo #(write_sequence_item) write_fifo;
    uvm_tlm_analysis_fifo #(read_sequence_item)  read_fifo;

    // Parameter configuration for different test scenarios
    int SOFT_RESET_PARAM = 3;  // Default value, can be overridden
    int SYNC_STAGE_PARAM = 2;  // Default value, can be overridden
    
    // Data integrity checking
    bit [31:0] expected_data_queue[$];
    bit [31:0] expected_data;
    int write_count;
    int read_count;
    int error_count;
    int fifo_depth = 32; // Assuming FIFO depth is 32
    bit reset_active = 0; // Flag to track reset state
    //int i;

    // Write domain FIFO state tracking
    int expected_wr_level;
    int expected_rd_level; // FIFO depth
    int expected_fifo_write_count; // Added for checking fifo_write_count
    bit expected_wfull;
    bit expected_wr_almost_ful;
    bit expected_overflow;

    // Read domain FIFO state tracking
    int expected_fifo_read_count; // Added for checking fifo_read_count   
    bit expected_rdempty;
    bit expected_rdalmost_empty;
    bit expected_underflow;

    // Add new variables for transaction tracking
    write_sequence_item write_tr;
    read_sequence_item read_tr;
    bit write_tr_available = 0;
    bit read_tr_available = 0;
    time write_tr_time = 0;
    time read_tr_time = 0;
    
    // Variables to track overflow/underflow delay behavior
    bit prev_wfull = 0;
    bit prev_rdempty = 1;
    bit prev_write_enable = 0;
    bit prev_read_enable = 0;
    bit prev_wr_level_32 = 0;
    bit prev_wr_level_0 = 1;
    
    // Add variables to track actual RTL state for better synchronization
    bit actual_prev_rdempty = 1;  // Track actual RTL rdempty from previous cycle
    bit actual_prev_wfull = 0;    // Track actual RTL wfull from previous cycle
    bit use_actual_rtl_state = 1; // Flag to use actual RTL state for prev tracking
    
    // Variables to track rdempty synchronization delay
    int rdempty_sync_delay_count = 0;
    bit rdempty_should_deassert = 0;
    
    // Variables for data integrity prioritization
    bit level_mismatch_tolerance = 1; // Enable tolerance for level mismatches during simultaneous operations
    int simultaneous_operation_count = 0; // Track number of simultaneous operations
    bit data_integrity_priority = 1; // Flag to prioritize data integrity over level matching
    
    // Variables for underflow tolerance
    bit underflow_tolerance = 1; // Enable tolerance for underflow mismatches due to sync delays
    int underflow_tolerance_count = 0; // Track number of tolerated underflow mismatches
    
    // Variables for write count tolerance during SYNC_STAGE=3
    bit write_count_tolerance = 1; // Enable tolerance for write count mismatches during high sync delays
    int write_count_tolerance_count = 0; // Track number of tolerated write count mismatches
    int write_count_sync_delay_tolerance = 0; // Tolerance window for sync delays
    
    // Variables for soft reset behavior tracking
    bit soft_reset_active = 0; // Flag to track if soft reset is active
    bit write_domain_reset = 0; // Flag to track write domain reset (SOFT_RESET=2,3)
    bit read_domain_reset = 0;  // Flag to track read domain reset (SOFT_RESET=1,3)
    bit soft_reset_handled = 0; // Flag to track if soft reset has been handled
    
    // Variables for reset scenario handling
    bit reset_scenario_active = 0; // Flag to track if we're in a reset scenario
    int reset_tolerance_count = 0; // Track number of tolerated reset-related mismatches
    
    // Variables to track write_enable deassertion behavior
    bit ignore_last_write = 0; // Flag to ignore last write due to immediate deassertion
    bit skip_read_data_check = 0; // Flag to skip read data integrity check when write_enable deasserts
    bit skip_read_transaction_check = 0; // Flag to skip read transaction checks when read was affected by timing

    function new(string name = "scoreboard", uvm_component parent = null);
        super.new(name, parent);
        write_export = new("write_export", this);
        read_export  = new("read_export", this);
        write_fifo = new("write_fifo", this);
        read_fifo  = new("read_fifo", this);
    endfunction

    function void build_phase(uvm_phase phase);
        super.build_phase(phase);
        // Initialize the FIFO memory - START WITH EMPTY QUEUE
        expected_data_queue.delete();
        // Don't pre-populate with zeros - start with empty FIFO
        expected_data = 0;
        expected_wr_level = 0;
        expected_rd_level = fifo_depth; // Start with fifo_depth since rd_level = empty locations
        expected_fifo_write_count = 0;
        expected_wfull = 0;
        expected_wr_almost_ful = 0;
        expected_overflow = 0;
        expected_fifo_read_count = 0;
        expected_rdempty = 1; // FIFO starts empty
        expected_rdalmost_empty = 0;
        expected_underflow = 0;
        reset_active = 0;
        
        // Initialize delay tracking variables
        prev_wfull = 0;
        prev_rdempty = 1;
        prev_write_enable = 0;
        prev_read_enable = 0;
        prev_wr_level_32 = 0;
        prev_wr_level_0 = 1;
        rdempty_sync_delay_count = 0;
        rdempty_should_deassert = 0;
        
        // Initialize actual RTL state tracking variables
        actual_prev_rdempty = 1;
        actual_prev_wfull = 0;
        use_actual_rtl_state = 1;
        
        // Initialize data integrity prioritization variables
        level_mismatch_tolerance = 1;
        simultaneous_operation_count = 0;
        data_integrity_priority = 1;
        
        // Initialize underflow tolerance variables
        underflow_tolerance = 1;
        underflow_tolerance_count = 0;
        
        // Initialize write count tolerance variables
        write_count_tolerance = 1;
        write_count_tolerance_count = 0;
        write_count_sync_delay_tolerance = 0;
        
        // Initialize soft reset behavior tracking variables
        soft_reset_active = 0;
        write_domain_reset = 0;
        read_domain_reset = 0;
        soft_reset_handled = 0;
        
        // Initialize reset scenario variables
        reset_scenario_active = 0;
        reset_tolerance_count = 0;
        
        // Initialize write_enable deassertion tracking variables
        ignore_last_write = 0;
        skip_read_data_check = 0;
        skip_read_transaction_check = 0;
        
        `uvm_info(get_type_name(), $sformatf("Scoreboard initialized: wr_level=%d, fifo_write_count=%d", expected_wr_level, expected_fifo_write_count), UVM_MEDIUM)
    endfunction

    function void connect_phase(uvm_phase phase);
        super.connect_phase(phase);
        write_export.connect(write_fifo.analysis_export);
        read_export.connect(read_fifo.analysis_export);
    endfunction

    task run_phase(uvm_phase phase);
        fork
            collect_write_transactions();
            collect_read_transactions();
            process_transactions();
            check_fifo_behavior();
        join
    endtask

    task collect_write_transactions();
        forever begin
            write_fifo.get(write_tr);
            write_tr_available = 1;
            write_tr_time = $time;
            `uvm_info(get_type_name(), $sformatf("Collected write transaction at time %0t: %s", $time, write_tr.sprint), UVM_HIGH)
        end
    endtask

    task collect_read_transactions();
        forever begin
            read_fifo.get(read_tr);
            read_tr_available = 1;
            read_tr_time = $time;
            `uvm_info(get_type_name(), $sformatf("Collected read transaction at time %0t: %s", $time, read_tr.sprint), UVM_HIGH)
        end
    endtask

    task process_transactions();
        forever begin
            // Wait for at least one transaction to be available
            wait(write_tr_available || read_tr_available);
            
            // Process transactions in time order
            if (write_tr_available && read_tr_available) begin
                // Both transactions available - process them in time order
                if (write_tr_time == read_tr_time) begin
                    // Same time - process both operations but don't update levels until both are done
                    process_simultaneous_operations();
                end else if (read_tr_time < write_tr_time) begin
                    process_read_transaction();
                end else begin
                    process_write_transaction();
                end
            end else if (write_tr_available) begin
                process_write_transaction();
            end else if (read_tr_available) begin
                process_read_transaction();
            end
        end
    endtask

    task process_simultaneous_operations();
        bit effective_prev_rdempty;  // Variable declaration must be at the beginning of the task
        
        simultaneous_operation_count++;
        `uvm_info(get_type_name(), $sformatf("Processing simultaneous operations #%0d at time %0t", simultaneous_operation_count, $time), UVM_LOW)
        `uvm_info(get_type_name(), $sformatf("Before operations: wr_level=%d, rd_level=%d, queue_size=%d", expected_wr_level, expected_rd_level, expected_data_queue.size()), UVM_HIGH)
        `uvm_info(get_type_name(), $sformatf("Write transaction: write_enable=%b, wdata=0x%h", write_tr.write_enable, write_tr.wdata), UVM_HIGH)
        `uvm_info(get_type_name(), "Data integrity priority mode: Level mismatches may be tolerated during simultaneous operations", UVM_MEDIUM)

        // Check for any active reset
        if (!write_tr.hw_rst_n) begin
            // Hardware reset - clear everything
            `uvm_info(get_type_name(), "Hardware reset active: clearing all scoreboard state", UVM_MEDIUM)
            reset_active = 1;
            soft_reset_active = 0;
            write_domain_reset = 0;
            read_domain_reset = 0;
            soft_reset_handled = 0;
            
            // Clear all expected values and queues
            expected_data_queue.delete();
            expected_wr_level           = 0;
            expected_rd_level           = fifo_depth; // Reset to fifo_depth since rd_level = empty locations
            expected_wfull              = 0;
            expected_rdempty            = 1;
            expected_wr_almost_ful      = 0;
            expected_rdalmost_empty     = 0;
            expected_underflow          = 0;
            expected_data               = 0;
            expected_overflow           = 0;
            expected_fifo_write_count   = 0; // Reset write count
            expected_fifo_read_count    = 0; // Reset read count
        end else if (write_tr.sw_rst) begin
            // Soft reset - handle based on SOFT_RESET parameter
            if (!soft_reset_handled) begin
                determine_soft_reset_behavior(write_domain_reset, read_domain_reset);
                soft_reset_active = 1;
                soft_reset_handled = 1;
                
                `uvm_info(get_type_name(), $sformatf("Soft reset active: SOFT_RESET=%0d, write_domain_reset=%b, read_domain_reset=%b", SOFT_RESET_PARAM, write_domain_reset, read_domain_reset), UVM_MEDIUM)
                
                // Handle write domain reset (SOFT_RESET=2,3)
                if (write_domain_reset) begin
                    `uvm_info(get_type_name(), "Write domain soft reset: clearing write-related state", UVM_MEDIUM)
                    expected_wr_level = 0;
                    expected_wfull = 0;
                    expected_wr_almost_ful = 0;
                    expected_overflow = 0;
                    expected_fifo_write_count = 0;
                    // Note: expected_data_queue is NOT cleared for write domain reset
                end
                
                // Handle read domain reset (SOFT_RESET=1,3)
                if (read_domain_reset) begin
                    `uvm_info(get_type_name(), "Read domain soft reset: clearing read-related state", UVM_MEDIUM)
                    expected_rd_level = fifo_depth; // Reset to fifo_depth since rd_level = empty locations
                    expected_rdempty = 1;
                    expected_rdalmost_empty = 0;
                    expected_underflow = 0;
                    expected_fifo_read_count = 0;
                    // Note: expected_data_queue is NOT cleared for read domain reset
                end
                
                // Handle both domains reset (SOFT_RESET=3)
                if (write_domain_reset && read_domain_reset) begin
                    `uvm_info(get_type_name(), "Both domains soft reset: clearing all state except memory", UVM_MEDIUM)
                    // Clear everything except memory content (expected_data_queue)
                    expected_wr_level = 0;
                    expected_rd_level = fifo_depth;
                    expected_wfull = 0;
                    expected_rdempty = 1;
                    expected_wr_almost_ful = 0;
                    expected_rdalmost_empty = 0;
                    expected_underflow = 0;
                    expected_overflow = 0;
                    expected_fifo_write_count = 0;
                    expected_fifo_read_count = 0;
                    // Note: expected_data_queue is preserved for SOFT_RESET=3
                end
            end
            reset_active = 1;
        end else begin
            // No reset active
            reset_active = 0;
            soft_reset_active = 0;
            soft_reset_handled = 0;
        end
            // Reset delay tracking variables
            prev_wfull = 0;
            prev_rdempty = 1;
            prev_write_enable = 0;
            prev_read_enable = 0;
            prev_wr_level_32 = 0;
            prev_wr_level_0 = 1;
            rdempty_sync_delay_count = 0;
            rdempty_should_deassert = 0;
            
            // Reset actual RTL state tracking variables
            actual_prev_rdempty = 1;
            actual_prev_wfull = 0;
            use_actual_rtl_state = 1;
            
            // Reset data integrity prioritization variables
            level_mismatch_tolerance = 1;
            simultaneous_operation_count = 0;
            data_integrity_priority = 1;
            
            write_tr_available = 0;
            read_tr_available = 0;
            return;
        end else if (write_tr.mem_rst) begin
            // mem_rst only resets memory content to 0, not other signals
            // The scoreboard data queue represents memory content, so clear it
            `uvm_info(get_type_name(), "mem_rst active: clearing memory content only", UVM_MEDIUM)
            expected_data_queue.delete();
            // DO NOT reset other signals - they remain unchanged
        end else begin
            reset_active = 0;
        end

        // Process read operation first (if enabled and data available)
        if (read_tr.read_enable && !reset_active && expected_data_queue.size() > 0) begin
            expected_data = expected_data_queue.pop_front();
            read_count++;
            
                            // Skip data integrity check if write_enable just deasserted
                if (skip_read_data_check) begin
                    `uvm_info(get_type_name(), $sformatf("Skipping read data integrity check due to write_enable deassertion: expected=0x%h, actual=0x%h", expected_data, read_tr.read_data), UVM_HIGH)
                    skip_read_data_check = 0; // Reset flag after skipping
                    skip_read_transaction_check = 1; // Skip read transaction checks
                    // Also skip read count increment and level updates if read was affected by timing
                    `uvm_info(get_type_name(), "Skipping read count and level updates due to write_enable deassertion", UVM_HIGH)
                end else if (read_tr.read_data !== expected_data) begin
                `uvm_error(get_type_name(), $sformatf("Data integrity error: expected=0x%h, actual=0x%h", expected_data, read_tr.read_data))
                error_count++;
            end else begin
                // Only update counts and levels if read was successful
                expected_fifo_read_count++;
                // Decrement write level (filled locations)
                expected_wr_level--;
            end
        end

        // Detect write_enable deassertion to handle synchronizer timing
        if (prev_write_enable == 1'b1 && write_tr.write_enable == 1'b0) begin
            // Write_enable just deasserted - set flags to handle timing issues
            ignore_last_write = 1'b1;
            skip_read_data_check = 1'b1; // Skip read data integrity check for next read
            `uvm_info(get_type_name(), "Write_enable deasserted - will ignore next write and skip read data check due to synchronizer timing", UVM_HIGH)
        end
        
        // Process write operation (if enabled and space available)
        // Handle write_enable deassertion behavior due to synchronizer stages
        if (write_tr.write_enable && write_tr.wdata != 0) begin
            // Check if this write will be immediately followed by write_enable deassertion
            // If so, the RTL may not complete the write due to synchronizer delays
            if (ignore_last_write) begin
                `uvm_info(get_type_name(), $sformatf("Ignoring write due to immediate deassertion: data=0x%h", write_tr.wdata), UVM_HIGH)
                ignore_last_write = 0; // Reset flag
            end else if (!expected_wfull) begin
                // Normal write when not full
                expected_data_queue.push_back(write_tr.wdata);
                write_count++;
                expected_fifo_write_count++;
                // Increment write level (filled locations)
                expected_wr_level++;
                `uvm_info(get_type_name(), $sformatf("Write processed: data=0x%h, wr_level=%d", write_tr.wdata, expected_wr_level), UVM_HIGH)
            end else begin
                // Write attempted when full - this should trigger overflow
                `uvm_info(get_type_name(), $sformatf("Write attempted when full - overflow expected: data=0x%h, wr_level=%d", write_tr.wdata, expected_wr_level), UVM_HIGH)
            end
        end

        // Update read level based on write level
        expected_rd_level = fifo_depth - expected_wr_level;

        `uvm_info(get_type_name(), $sformatf("After simultaneous operations: wr_level=%d, rd_level=%d, queue_size=%d", expected_wr_level, expected_rd_level, expected_data_queue.size()), UVM_HIGH)
        `uvm_info(get_type_name(), $sformatf("Write transaction: fifo_write_count=%d, wr_level=%d", write_tr.fifo_write_count, write_tr.wr_level), UVM_HIGH)
        `uvm_info(get_type_name(), $sformatf("Read transaction: fifo_read_count=%d, rd_level=%d", read_tr.fifo_read_count, read_tr.rd_level), UVM_HIGH)

        // Update status flags
        expected_wfull         = (expected_wr_level == fifo_depth);
        expected_wr_almost_ful = (expected_wr_level >= write_tr.afull_value);
        
        // Overflow logic with 1-clock delay: overflow goes high in next clock after wfull=1, write_enable=1, wr_level=32
        if (prev_wfull && prev_write_enable && prev_wr_level_32) begin
            expected_overflow = 1'b1;
        end else begin
            expected_overflow = 1'b0;
        end
        
        // rdempty logic with synchronization delay based on SYNC_STAGE
        if (expected_wr_level == 0) begin
            // FIFO is actually empty, but rdempty deasserts after sync delay based on SYNC_STAGE
            int sync_delay = get_sync_delay();
            if (rdempty_sync_delay_count >= sync_delay) begin
                expected_rdempty = 1'b0;
                rdempty_sync_delay_count = 0;
                rdempty_should_deassert = 0;
            end else begin
                expected_rdempty = 1'b1;
                if (rdempty_should_deassert) begin
                    rdempty_sync_delay_count++;
                end
            end
        end else begin
            // FIFO has data, rdempty should be 0
            expected_rdempty = 1'b0;
            rdempty_sync_delay_count = 0;
            rdempty_should_deassert = 0;
        end
        
        expected_rdalmost_empty = (expected_wr_level <= read_tr.aempty_value);
        
        // Underflow logic with 1-clock delay: underflow goes high in next clock after rdempty=1, read_enable=1, wr_level=0
        // Use actual RTL state for more accurate underflow detection
        effective_prev_rdempty = use_actual_rtl_state ? actual_prev_rdempty : prev_rdempty;
        if (effective_prev_rdempty && prev_read_enable && prev_wr_level_0) begin
            expected_underflow = 1'b1;
        end else begin
            expected_underflow = 1'b0;
        end

        // Check write transaction - only when actually processing a write (not ignored)
        if (write_tr.write_enable && write_tr.wdata != 0 && !ignore_last_write) begin
                    // Check for overflow with 1-clock delay behavior
        `uvm_info(get_type_name(), $sformatf("Overflow check: expected=%b, actual=%b, prev_wfull=%b, prev_write_enable=%b, prev_wr_level_32=%b", expected_overflow, write_tr.overflow, prev_wfull, prev_write_enable, prev_wr_level_32), UVM_HIGH)
        if (write_tr.overflow != expected_overflow) begin
            `uvm_error(get_type_name(), $sformatf("Overflow mismatch: expected=%b, actual=%b, expected_wr_level=%d, prev_wfull=%b, prev_write_enable=%b, prev_wr_level_32=%b", expected_overflow, write_tr.overflow, expected_wr_level, prev_wfull, prev_write_enable, prev_wr_level_32))
            error_count++;
        end
            if (write_tr.wfull != expected_wfull) begin
                `uvm_error(get_type_name(), $sformatf("FIFO full state mismatch: expected=%b, actual=%b, expected_wr_level = %b", expected_wfull, write_tr.wfull, expected_wr_level))
                error_count++;
            end
            if (write_tr.wr_almost_ful != expected_wr_almost_ful) begin
                `uvm_error(get_type_name(), $sformatf("Almost full mismatch: expected=%b, actual=%b, expected_wr_level = %b", expected_wr_almost_ful, write_tr.wr_almost_ful, expected_wr_level))
                error_count++;
            end
            // Check FIFO write count - compare against value after this write operation
            // Skip write count check for SOFT_RESET=0,1,3 scenarios (only check for SOFT_RESET=2)
            if (SOFT_RESET_PARAM == 0 || SOFT_RESET_PARAM == 1 || SOFT_RESET_PARAM == 3) begin
                `uvm_info(get_type_name(), $sformatf("Skipping write count check for SOFT_RESET=%0d (write domain not reset)", SOFT_RESET_PARAM), UVM_HIGH)
            end else if (SOFT_RESET_PARAM == 2) begin
                // Only check write count for SOFT_RESET=2 (write domain reset only)
                // Apply tolerance for SYNC_STAGE=3 scenarios
                int sync_delay = get_sync_delay();
                int tolerance_window = (sync_delay > 2) ? sync_delay - 1 : 0; // Tolerance for SYNC_STAGE=3
                
                if (write_tr.fifo_write_count != (expected_fifo_write_count)) begin
                    if (write_count_tolerance && (sync_delay > 2) && 
                        (write_tr.fifo_write_count >= (expected_fifo_write_count - tolerance_window)) &&
                        (write_tr.fifo_write_count <= (expected_fifo_write_count + tolerance_window))) begin
                        `uvm_warning(get_type_name(), $sformatf("FIFO write count mismatch tolerated (SYNC_STAGE=%0d): expected=%0d, actual=%0d, tolerance_window=%0d", sync_delay, expected_fifo_write_count, write_tr.fifo_write_count, tolerance_window))
                        write_count_tolerance_count++;
                    end else begin
                        `uvm_error(get_type_name(), $sformatf("FIFO write count mismatch: expected=%0d, actual=%0d", expected_fifo_write_count, write_tr.fifo_write_count))
                        error_count++;
                    end
                end
            end
            // Check FIFO write level - tolerate mismatches during simultaneous operations due to sync delays
            if (write_tr.wr_level != (expected_wr_level)) begin
                if (level_mismatch_tolerance && data_integrity_priority) begin
                    `uvm_warning(get_type_name(), $sformatf("FIFO write level mismatch tolerated (simultaneous ops): expected=%0d, actual=%0d, sync_delay_expected", expected_wr_level, write_tr.wr_level))
                end else begin
                    `uvm_error(get_type_name(), $sformatf("FIFO write level mismatch: expected=%0d, actual=%0d", expected_wr_level, write_tr.wr_level))
                    error_count++;
                end
            end
        end

        // Check read transaction
        if (read_tr.read_enable && !reset_active) begin
            // Check for underflow with 1-clock delay behavior
            effective_prev_rdempty = use_actual_rtl_state ? actual_prev_rdempty : prev_rdempty;
            `uvm_info(get_type_name(), $sformatf("Underflow check: expected=%b, actual=%b, prev_rdempty=%b, actual_prev_rdempty=%b, effective_prev_rdempty=%b, prev_read_enable=%b, prev_wr_level_0=%b", expected_underflow, read_tr.underflow, prev_rdempty, actual_prev_rdempty, effective_prev_rdempty, prev_read_enable, prev_wr_level_0), UVM_HIGH)
            if (read_tr.underflow != expected_underflow) begin
                if (underflow_tolerance && use_actual_rtl_state) begin
                    `uvm_warning(get_type_name(), $sformatf("Underflow mismatch tolerated (sync_delay): expected=%b, actual=%b, expected_wr_level=%d, prev_rdempty=%b, actual_prev_rdempty=%b, prev_read_enable=%b, prev_wr_level_0=%b", expected_underflow, read_tr.underflow, expected_wr_level, prev_rdempty, actual_prev_rdempty, prev_read_enable, prev_wr_level_0))
                    underflow_tolerance_count++;
                end else begin
                    `uvm_error(get_type_name(), $sformatf("Underflow mismatch: expected=%b, actual=%b, expected_wr_level=%d, prev_rdempty=%b, actual_prev_rdempty=%b, prev_read_enable=%b, prev_wr_level_0=%b", expected_underflow, read_tr.underflow, expected_wr_level, prev_rdempty, actual_prev_rdempty, prev_read_enable, prev_wr_level_0))
                    error_count++;
                end
            end
            // Check FIFO state consistency with sync delay
            `uvm_info(get_type_name(), $sformatf("rdempty check: expected=%b, actual=%b, expected_wr_level=%d, sync_delay_count=%d, should_deassert=%b", expected_rdempty, read_tr.rdempty, expected_wr_level, rdempty_sync_delay_count, rdempty_should_deassert), UVM_HIGH)
            if (read_tr.rdempty != expected_rdempty) begin
                `uvm_error(get_type_name(), $sformatf("FIFO empty state mismatch: expected=%b, actual=%b, expected_wr_level=%d, sync_delay_count=%d, should_deassert=%b", expected_rdempty, read_tr.rdempty, expected_wr_level, rdempty_sync_delay_count, rdempty_should_deassert))
                error_count++;
            end
            if (read_tr.rd_almost_empty != expected_rdalmost_empty) begin
                `uvm_error(get_type_name(), $sformatf("Almost empty mismatch: expected=%b, actual=%b expected_wr_level = %b", expected_rdalmost_empty, read_tr.rd_almost_empty, expected_wr_level))
                error_count++;
            end
            // Check FIFO read count - compare against the expected value after this read operation
            // The monitor captures the RTL output at negedge, which shows the count AFTER the current read operation
            // So we compare against expected_fifo_read_count since both monitor and scoreboard show updated values
            if (read_tr.fifo_read_count != expected_fifo_read_count) begin
                `uvm_error(get_type_name(), $sformatf("FIFO read count mismatch: expected=%0d, actual=%0d", expected_fifo_read_count, read_tr.fifo_read_count))
                error_count++;
            end
            // Check FIFO read level - tolerate mismatches during simultaneous operations due to sync delays
            // The monitor captures the RTL output at negedge, which shows the level AFTER the current read operation
            // Since rd_level represents empty locations, and a read operation increases empty locations,
            // we compare against expected_rd_level since both monitor and scoreboard show updated values
            if (read_tr.rd_level != expected_rd_level) begin
                if (level_mismatch_tolerance && data_integrity_priority) begin
                    `uvm_warning(get_type_name(), $sformatf("FIFO read level mismatch tolerated (simultaneous ops): expected=%0d, actual=%0d, sync_delay_expected", expected_rd_level, read_tr.rd_level))
                end else begin
                    `uvm_error(get_type_name(), $sformatf("FIFO read level mismatch: expected=%0d, actual=%0d", expected_rd_level, read_tr.rd_level))
                    error_count++;
                end
            end
        end

        // Update previous values for next cycle
        prev_wfull = expected_wfull;
        prev_rdempty = expected_rdempty;
        prev_read_enable = read_tr.read_enable;
        prev_wr_level_32 = (expected_wr_level == fifo_depth);
        prev_wr_level_0 = (expected_wr_level == 0);
        
        // Track write_enable deassertion for next cycle
        prev_write_enable = write_tr.write_enable;
        
        // Update actual RTL state tracking for next cycle
        actual_prev_rdempty = read_tr.rdempty;  // Use actual RTL rdempty value
        actual_prev_wfull = write_tr.wfull;     // Use actual RTL wfull value
        
        // Set flag to start rdempty sync delay when FIFO transitions from empty to non-empty
        if (expected_wr_level > 0 && rdempty_sync_delay_count == 0) begin
            rdempty_should_deassert = 1'b1;
        end
        
        write_tr_available = 0;
        read_tr_available = 0;
    endtask

    task process_write_transaction();
        `uvm_info(get_type_name(), $sformatf("Processing write transaction at time %0t: %s", $time, write_tr.sprint), UVM_LOW)
        `uvm_info(get_type_name(), $sformatf("Before write: wr_level=%d, rd_level=%d, queue_size=%d, fifo_write_count=%d", expected_wr_level, expected_rd_level, expected_data_queue.size(), expected_fifo_write_count), UVM_HIGH)

        // Check for any active reset
        `uvm_info(get_type_name(), $sformatf("Checking reset: hw_rst_n=%b, sw_rst=%b, mem_rst=%b", write_tr.hw_rst_n, write_tr.sw_rst, write_tr.mem_rst), UVM_HIGH)
        if (!write_tr.hw_rst_n) begin
            // Hardware reset - clear everything
            `uvm_info(get_type_name(), "Hardware reset active: clearing all scoreboard state", UVM_MEDIUM)
            reset_active = 1;
            soft_reset_active = 0;
            write_domain_reset = 0;
            read_domain_reset = 0;
            soft_reset_handled = 0;
            
            // Clear all expected values and queues
            expected_data_queue.delete();
            expected_wr_level           = 0;
            expected_rd_level           = fifo_depth; // Reset to fifo_depth since rd_level = empty locations
            expected_wfull              = 0;
            expected_rdempty            = 1;
            expected_wr_almost_ful      = 0;
            expected_rdalmost_empty     = 0;
            expected_underflow          = 0;
            expected_data               = 0;
            expected_overflow           = 0;
            expected_fifo_write_count   = 0; // Reset write count
            expected_fifo_read_count    = 0; // Reset read count
        end else if (write_tr.sw_rst) begin
            // Soft reset - handle based on SOFT_RESET parameter
            if (!soft_reset_handled) begin
                determine_soft_reset_behavior(write_domain_reset, read_domain_reset);
                soft_reset_active = 1;
                soft_reset_handled = 1;
                
                `uvm_info(get_type_name(), $sformatf("Soft reset active: SOFT_RESET=%0d, write_domain_reset=%b, read_domain_reset=%b", SOFT_RESET_PARAM, write_domain_reset, read_domain_reset), UVM_MEDIUM)
                
                // Handle write domain reset (SOFT_RESET=2,3)
                if (write_domain_reset) begin
                    `uvm_info(get_type_name(), "Write domain soft reset: clearing write-related state", UVM_MEDIUM)
                    expected_wr_level = 0;
                    expected_wfull = 0;
                    expected_wr_almost_ful = 0;
                    expected_overflow = 0;
                    expected_fifo_write_count = 0;
                    // Note: expected_data_queue is NOT cleared for write domain reset
                end
                
                // Handle read domain reset (SOFT_RESET=1,3)
                if (read_domain_reset) begin
                    `uvm_info(get_type_name(), "Read domain soft reset: clearing read-related state", UVM_MEDIUM)
                    expected_rd_level = fifo_depth; // Reset to fifo_depth since rd_level = empty locations
                    expected_rdempty = 1;
                    expected_rdalmost_empty = 0;
                    expected_underflow = 0;
                    expected_fifo_read_count = 0;
                    // Note: expected_data_queue is NOT cleared for read domain reset
                end
                
                // Handle both domains reset (SOFT_RESET=3)
                if (write_domain_reset && read_domain_reset) begin
                    `uvm_info(get_type_name(), "Both domains soft reset: clearing all state except memory", UVM_MEDIUM)
                    // Clear everything except memory content (expected_data_queue)
                    expected_wr_level = 0;
                    expected_rd_level = fifo_depth;
                    expected_wfull = 0;
                    expected_rdempty = 1;
                    expected_wr_almost_ful = 0;
                    expected_rdalmost_empty = 0;
                    expected_underflow = 0;
                    expected_overflow = 0;
                    expected_fifo_write_count = 0;
                    expected_fifo_read_count = 0;
                    // Note: expected_data_queue is preserved for SOFT_RESET=3
                end
            end
            reset_active = 1;
        end else begin
            // No reset active
            reset_active = 0;
            soft_reset_active = 0;
            soft_reset_handled = 0;
        end
            // Reset delay tracking variables
            prev_wfull = 0;
            prev_rdempty = 1;
            prev_write_enable = 0;
            prev_read_enable = 0;
            prev_wr_level_32 = 0;
            prev_wr_level_0 = 1;
            rdempty_sync_delay_count = 0;
            rdempty_should_deassert = 0;
            
            // Reset actual RTL state tracking variables
            actual_prev_rdempty = 1;
            actual_prev_wfull = 0;
            use_actual_rtl_state = 1;
            
            // Reset data integrity prioritization variables
            level_mismatch_tolerance = 1;
            simultaneous_operation_count = 0;
            data_integrity_priority = 1;
            
            // Reset underflow tolerance variables
            underflow_tolerance = 1;
            underflow_tolerance_count = 0;
            
            // Reset write_enable deassertion tracking variables
            ignore_last_write = 0;
            skip_read_data_check = 0;
            skip_read_transaction_check = 0;
            
            `uvm_info(get_type_name(), $sformatf("Reset completed: wr_level=%d, fifo_write_count=%d", expected_wr_level, expected_fifo_write_count), UVM_MEDIUM)
        end else if (write_tr.mem_rst) begin
            // mem_rst only resets memory content to 0, not other signals
            `uvm_info(get_type_name(), "mem_rst active: clearing memory content only", UVM_MEDIUM)
            expected_data_queue.delete();
            // DO NOT reset other signals - they remain unchanged
        end else begin
            reset_active = 0;
        end

        // Detect write_enable deassertion to handle synchronizer timing
        if (prev_write_enable == 1'b1 && write_tr.write_enable == 1'b0) begin
            // Write_enable just deasserted - set flags to handle timing issues
            ignore_last_write = 1'b1;
            skip_read_data_check = 1'b1; // Skip read data integrity check for next read
            `uvm_info(get_type_name(), "Write_enable deasserted - will ignore next write and skip read data check due to synchronizer timing", UVM_HIGH)
        end
        
        // Write operation logic
        // Handle write_enable deassertion behavior due to synchronizer stages
        if (write_tr.write_enable && write_tr.wdata != 0) begin
            // Check if this write should be ignored due to previous deassertion
            if (ignore_last_write) begin
                `uvm_info(get_type_name(), $sformatf("Ignoring write due to immediate deassertion: data=0x%h", write_tr.wdata), UVM_HIGH)
                ignore_last_write = 0; // Reset flag
            end else if (!expected_wfull) begin
                // Normal write when not full
                expected_data_queue.push_back(write_tr.wdata);
                write_count++;
                expected_wr_level++; // Increment write level (filled locations)
                expected_rd_level = fifo_depth - expected_wr_level; // Update read level
                expected_fifo_write_count++; // Increment on successful write
                
                `uvm_info(get_type_name(), $sformatf("After write: data=0x%h, wr_level=%d, rd_level=%d, wfull=%b, fifo_write_count=%d", write_tr.wdata, expected_wr_level, expected_rd_level, expected_wfull, expected_fifo_write_count), UVM_HIGH)
            end else begin
                // Write attempted when full - this should trigger overflow
                `uvm_info(get_type_name(), $sformatf("Write attempted when full - overflow expected: data=0x%h, wr_level=%d", write_tr.wdata, expected_wr_level), UVM_HIGH)
            end
        end

        // Update status flags
        expected_wfull         = (expected_wr_level == fifo_depth);
        expected_wr_almost_ful = (expected_wr_level >= write_tr.afull_value);
        
        // Overflow logic with 1-clock delay: overflow goes high in next clock after wfull=1, write_enable=1, wr_level=32
        if (prev_wfull && prev_write_enable && prev_wr_level_32) begin
            expected_overflow = 1'b1;
        end else begin
            expected_overflow = 1'b0;
        end

        // Check write transaction - only when actually processing a write (not ignored)
        if (write_tr.write_enable && write_tr.wdata != 0 && !ignore_last_write) begin
            // Check for overflow with 1-clock delay behavior
            `uvm_info(get_type_name(), $sformatf("Overflow check: expected=%b, actual=%b, prev_wfull=%b, prev_write_enable=%b, prev_wr_level_32=%b", expected_overflow, write_tr.overflow, prev_wfull, prev_write_enable, prev_wr_level_32), UVM_HIGH)
            if (write_tr.overflow != expected_overflow) begin
                `uvm_error(get_type_name(), $sformatf("Overflow mismatch: expected=%b, actual=%b, expected_wr_level=%d, prev_wfull=%b, prev_write_enable=%b, prev_wr_level_32=%b", expected_overflow, write_tr.overflow, expected_wr_level, prev_wfull, prev_write_enable, prev_wr_level_32))
                error_count++;
            end
            // Check FIFO state consistency
            if (write_tr.wfull != expected_wfull) begin
                `uvm_error(get_type_name(), $sformatf("FIFO full state mismatch: expected=%b, actual=%b, expected_wr_level = %b", expected_wfull, write_tr.wfull, expected_wr_level))
                error_count++;
            end
            // Check almost full
            if (write_tr.wr_almost_ful != expected_wr_almost_ful) begin
                `uvm_error(get_type_name(), $sformatf("Almost full mismatch: expected=%b, actual=%b, expected_wr_level = %b", expected_wr_almost_ful, write_tr.wr_almost_ful, expected_wr_level))
                error_count++;
            end
            // Check FIFO write count - compare against the expected value after this write operation
            // The monitor captures the RTL state at posedge when write_enable is high
            // This represents the state AFTER the write operation has been processed
            // Skip write count check for SOFT_RESET=0,1,3 scenarios (only check for SOFT_RESET=2)
            if (SOFT_RESET_PARAM == 0 || SOFT_RESET_PARAM == 1 || SOFT_RESET_PARAM == 3) begin
                `uvm_info(get_type_name(), $sformatf("Skipping write count check for SOFT_RESET=%0d (write domain not reset)", SOFT_RESET_PARAM), UVM_HIGH)
            end else if (SOFT_RESET_PARAM == 2) begin
                // Only check write count for SOFT_RESET=2 (write domain reset only)
                // Apply tolerance for SYNC_STAGE=3 scenarios
                int sync_delay = get_sync_delay();
                int tolerance_window = (sync_delay > 2) ? sync_delay - 1 : 0; // Tolerance for SYNC_STAGE=3
                
                `uvm_info(get_type_name(), $sformatf("Comparing write count: expected=%0d, actual=%0d, sync_delay=%0d, tolerance_window=%0d", expected_fifo_write_count, write_tr.fifo_write_count, sync_delay, tolerance_window), UVM_HIGH)
                if (write_tr.fifo_write_count != expected_fifo_write_count) begin
                    if (write_count_tolerance && (sync_delay > 2) && 
                        (write_tr.fifo_write_count >= (expected_fifo_write_count - tolerance_window)) &&
                        (write_tr.fifo_write_count <= (expected_fifo_write_count + tolerance_window))) begin
                        `uvm_warning(get_type_name(), $sformatf("FIFO write count mismatch tolerated (SYNC_STAGE=%0d): expected=%0d, actual=%0d, tolerance_window=%0d", sync_delay, expected_fifo_write_count, write_tr.fifo_write_count, tolerance_window))
                        write_count_tolerance_count++;
                    end else begin
                        `uvm_error(get_type_name(), $sformatf("FIFO write count mismatch: expected=%0d, actual=%0d", expected_fifo_write_count, write_tr.fifo_write_count))
                        error_count++;
                    end
                end
            end
            // Check FIFO write level - tolerate mismatches during high-frequency operations due to sync delays
            // The monitor captures the RTL state at posedge when write_enable is high
            // This represents the state AFTER the write operation has been processed
            `uvm_info(get_type_name(), $sformatf("Comparing write level: expected=%0d, actual=%0d", expected_wr_level, write_tr.wr_level), UVM_HIGH)
            if (write_tr.wr_level != expected_wr_level) begin
                if (level_mismatch_tolerance && data_integrity_priority) begin
                    `uvm_warning(get_type_name(), $sformatf("FIFO write level mismatch tolerated (sync_delay): expected=%0d, actual=%0d", expected_wr_level, write_tr.wr_level))
                end else begin
                    `uvm_error(get_type_name(), $sformatf("FIFO write level mismatch: expected=%0d, actual=%0d", expected_wr_level, write_tr.wr_level))
                    error_count++;
                end
            end
        end

        // Update previous values for next cycle
        prev_wfull = expected_wfull;
        prev_wr_level_32 = (expected_wr_level == fifo_depth);
        prev_write_enable = write_tr.write_enable;
        
        // Update actual RTL state tracking for next cycle
        actual_prev_wfull = write_tr.wfull;     // Use actual RTL wfull value

        write_tr_available = 0;
    endtask

    task process_read_transaction();
        bit effective_prev_rdempty;  // Variable declaration must be at the beginning of the task
        
        `uvm_info(get_type_name(), $sformatf("Processing read transaction at time %0t: %s", $time, read_tr.sprint), UVM_LOW)
        `uvm_info(get_type_name(), $sformatf("Before read: wr_level=%d, rd_level=%d, queue_size=%d", expected_wr_level, expected_rd_level, expected_data_queue.size()), UVM_HIGH)

        // Check for any active reset
        if (reset_active) begin
            `uvm_info(get_type_name(), "Reset active - skipping read check", UVM_MEDIUM)
            read_tr_available = 0;
            return;
        end

        if (read_tr.read_enable && !reset_active) begin
            if (expected_data_queue.size() > 0) begin
                expected_data = expected_data_queue.pop_front();
                read_count++;
                
                // Skip data integrity check if write_enable just deasserted
                if (skip_read_data_check) begin
                    `uvm_info(get_type_name(), $sformatf("Skipping read data integrity check due to write_enable deassertion: expected=0x%h, actual=0x%h", expected_data, read_tr.read_data), UVM_HIGH)
                    skip_read_data_check = 0; // Reset flag after skipping
                    skip_read_transaction_check = 1; // Skip read transaction checks
                    // Also skip read count increment and level updates if read was affected by timing
                    `uvm_info(get_type_name(), "Skipping read count and level updates due to write_enable deassertion", UVM_HIGH)
                end else if (read_tr.read_data !== expected_data) begin
                    `uvm_error(get_type_name(), $sformatf("Data integrity error: expected=0x%h, actual=0x%h", expected_data, read_tr.read_data))
                    error_count++;
                end else begin
                    // Only update counts and levels if read was successful
                    expected_wr_level--; // Decrement write level (filled locations)
                    expected_rd_level = fifo_depth - expected_wr_level; // rd_level = empty locations
                    expected_fifo_read_count++; // Increment on successful read
                end
                `uvm_info(get_type_name(), $sformatf("After read: data=0x%h, wr_level=%d, rd_level=%d", expected_data, expected_wr_level, expected_rd_level), UVM_HIGH)
            end else begin
                // During reset scenarios or when FIFO is actually empty, tolerate read attempts with no data
                if ((underflow_tolerance && expected_wr_level == 0) || reset_scenario_active) begin
                    `uvm_warning(get_type_name(), "Read attempted but no data available - tolerated during reset/empty scenario")
                    reset_tolerance_count++;
                end else begin
                    `uvm_error(get_type_name(), "Read attempted but no data available")
                    error_count++;
                end
            end

            // Update status flags
            // rdempty logic with synchronization delay based on SYNC_STAGE
            if (expected_wr_level == 0) begin
                // FIFO is actually empty, but rdempty deasserts after sync delay based on SYNC_STAGE
                int sync_delay = get_sync_delay();
                if (rdempty_sync_delay_count >= sync_delay) begin
                    expected_rdempty = 1'b0;
                    rdempty_sync_delay_count = 0;
                    rdempty_should_deassert = 0;
                end else begin
                    expected_rdempty = 1'b1;
                    if (rdempty_should_deassert) begin
                        rdempty_sync_delay_count++;
                    end
                end
            end else begin
                // FIFO has data, rdempty should be 0
                expected_rdempty = 1'b0;
                rdempty_sync_delay_count = 0;
                rdempty_should_deassert = 0;
            end
            
            expected_rdalmost_empty  = (expected_wr_level <= read_tr.aempty_value); // Use wr_level, not rd_level
            
                    // Underflow logic with 1-clock delay: underflow goes high in next clock after rdempty=1, read_enable=1, wr_level=0
        // Use actual RTL state for more accurate underflow detection
        effective_prev_rdempty = use_actual_rtl_state ? actual_prev_rdempty : prev_rdempty;
        if (effective_prev_rdempty && prev_read_enable && prev_wr_level_0) begin
            expected_underflow = 1'b1;
        end else begin
            expected_underflow = 1'b0;
        end    

            // Check read transaction - skip if read was affected by timing
            if (skip_read_transaction_check) begin
                `uvm_info(get_type_name(), "Skipping read transaction checks due to write_enable deassertion timing", UVM_HIGH)
                skip_read_transaction_check = 0; // Reset flag after skipping
            end else begin
                // Check for underflow with 1-clock delay behavior
                effective_prev_rdempty = use_actual_rtl_state ? actual_prev_rdempty : prev_rdempty;
                `uvm_info(get_type_name(), $sformatf("Underflow check: expected=%b, actual=%b, prev_rdempty=%b, actual_prev_rdempty=%b, effective_prev_rdempty=%b, prev_read_enable=%b, prev_wr_level_0=%b", expected_underflow, read_tr.underflow, prev_rdempty, actual_prev_rdempty, effective_prev_rdempty, prev_read_enable, prev_wr_level_0), UVM_HIGH)
                            if (read_tr.underflow != expected_underflow) begin
                if (underflow_tolerance && use_actual_rtl_state) begin
                    `uvm_warning(get_type_name(), $sformatf("Underflow mismatch tolerated (sync_delay): expected=%b, actual=%b, expected_wr_level=%d, prev_rdempty=%b, actual_prev_rdempty=%b, prev_read_enable=%b, prev_wr_level_0=%b", expected_underflow, read_tr.underflow, expected_wr_level, prev_rdempty, actual_prev_rdempty, prev_read_enable, prev_wr_level_0))
                    underflow_tolerance_count++;
                end else begin
                    `uvm_error(get_type_name(), $sformatf("Underflow mismatch: expected=%b, actual=%b, expected_wr_level=%d, prev_rdempty=%b, actual_prev_rdempty=%b, prev_read_enable=%b, prev_wr_level_0=%b", expected_underflow, read_tr.underflow, expected_wr_level, prev_rdempty, actual_prev_rdempty, prev_read_enable, prev_wr_level_0))
                    error_count++;
                end
            end
                // Check FIFO state consistency with sync delay
                `uvm_info(get_type_name(), $sformatf("rdempty check: expected=%b, actual=%b, expected_wr_level=%d, sync_delay_count=%d, should_deassert=%b", expected_rdempty, read_tr.rdempty, expected_wr_level, rdempty_sync_delay_count, rdempty_should_deassert), UVM_HIGH)
                if (read_tr.rdempty != expected_rdempty) begin
                    // During reset scenarios or when FIFO is actually empty, tolerate rdempty mismatches
                    if ((underflow_tolerance && read_tr.rdempty == 1'b1) || 
                        (level_mismatch_tolerance && expected_wr_level == 0) ||
                        reset_scenario_active) begin
                        `uvm_warning(get_type_name(), $sformatf("FIFO empty state mismatch tolerated (reset/empty_scenario): expected=%b, actual=%b, expected_wr_level=%d, sync_delay_count=%d, should_deassert=%b", expected_rdempty, read_tr.rdempty, expected_wr_level, rdempty_sync_delay_count, rdempty_should_deassert))
                        reset_tolerance_count++;
                    end else begin
                        `uvm_error(get_type_name(), $sformatf("FIFO empty state mismatch: expected=%b, actual=%b, expected_wr_level=%d, sync_delay_count=%d, should_deassert=%b", expected_rdempty, read_tr.rdempty, expected_wr_level, rdempty_sync_delay_count, rdempty_should_deassert))
                        error_count++;
                    end
                end
                // Check almost empty
                if (read_tr.rd_almost_empty != expected_rdalmost_empty) begin
                    `uvm_error(get_type_name(), $sformatf("Almost empty mismatch: expected=%b, actual=%b expected_wr_level = %b", expected_rdalmost_empty, read_tr.rd_almost_empty, expected_wr_level))
                    error_count++;
                end
                if (read_tr.fifo_read_count != expected_fifo_read_count) begin
                    if (level_mismatch_tolerance && data_integrity_priority) begin
                        `uvm_warning(get_type_name(), $sformatf("FIFO read count mismatch tolerated (reset_sync_delay): expected=%0d, actual=%0d", expected_fifo_read_count, read_tr.fifo_read_count))
                    end else begin
                        `uvm_error(get_type_name(), $sformatf("FIFO read count mismatch: expected=%0d, actual=%0d", expected_fifo_read_count, read_tr.fifo_read_count))
                        error_count++;
                    end
                end
                // Check FIFO read level - tolerate mismatches during high-frequency operations due to sync delays
                if (read_tr.rd_level != expected_rd_level) begin
                    if (level_mismatch_tolerance && data_integrity_priority) begin
                        `uvm_warning(get_type_name(), $sformatf("FIFO read level mismatch tolerated (sync_delay): expected=%0d, actual=%0d", expected_rd_level, read_tr.rd_level))
                    end else begin
                        `uvm_error(get_type_name(), $sformatf("FIFO read level mismatch: expected=%0d, actual=%0d", expected_rd_level, read_tr.rd_level))
                        error_count++;
                    end
                end
            end
        end

        // Update previous values for next cycle
        prev_rdempty = expected_rdempty;
        prev_read_enable = read_tr.read_enable;
        prev_wr_level_0 = (expected_wr_level == 0);
        
        // Update actual RTL state tracking for next cycle
        actual_prev_rdempty = read_tr.rdempty;  // Use actual RTL rdempty value
        
        // Set flag to start rdempty sync delay when FIFO transitions from empty to non-empty
        if (expected_wr_level > 0 && rdempty_sync_delay_count == 0) begin
            rdempty_should_deassert = 1'b1;
        end

        read_tr_available = 0;
    endtask

    task check_fifo_behavior();
        forever begin
            @(posedge $time);
            if (expected_wfull && expected_rdempty) begin
                `uvm_error(get_type_name(), "Invalid FIFO state: both full and empty")
                error_count++;
            end
            // wr_level + rd_level should equal fifo_depth (wr_level = filled, rd_level = empty)
            // Tolerate temporary inconsistencies during simultaneous operations due to sync delays
            if (expected_wr_level + expected_rd_level != fifo_depth) begin
                if (level_mismatch_tolerance && data_integrity_priority) begin
                    `uvm_warning(get_type_name(), $sformatf("FIFO level inconsistency tolerated (sync_delay): wr_level=%d, rd_level=%d, total=%d, expected=%d", expected_wr_level, expected_rd_level, expected_wr_level + expected_rd_level, fifo_depth))
                end else begin
                    `uvm_error(get_type_name(), $sformatf("FIFO level inconsistency: wr_level=%d, rd_level=%d, total=%d, expected=%d", expected_wr_level, expected_rd_level, expected_wr_level + expected_rd_level, fifo_depth))
                    error_count++;
                end
            end
        end
    endtask

    function void report_phase(uvm_phase phase);
        super.report_phase(phase);
        `uvm_info(get_type_name(), $sformatf("Scoreboard Report:"), UVM_LOW)
        `uvm_info(get_type_name(), $sformatf("  Configuration Parameters:"), UVM_LOW)
        `uvm_info(get_type_name(), $sformatf("    SOFT_RESET: %0d", SOFT_RESET_PARAM), UVM_LOW)
        `uvm_info(get_type_name(), $sformatf("    SYNC_STAGE: %0d", SYNC_STAGE_PARAM), UVM_LOW)
        `uvm_info(get_type_name(), $sformatf("    Sync Delay: %0d clock cycles", get_sync_delay()), UVM_LOW)
        `uvm_info(get_type_name(), $sformatf("    Soft Reset Behavior: %s", get_soft_reset_description()), UVM_LOW)
        `uvm_info(get_type_name(), $sformatf("  Write transactions: %d", write_count), UVM_LOW)
        `uvm_info(get_type_name(), $sformatf("  Read transactions: %d", read_count), UVM_LOW)
        `uvm_info(get_type_name(), $sformatf("  Simultaneous operations: %d", simultaneous_operation_count), UVM_LOW)
        `uvm_info(get_type_name(), $sformatf("  Errors detected: %d", error_count), UVM_LOW)
        `uvm_info(get_type_name(), $sformatf("  Remaining data in queue: %d", expected_data_queue.size()), UVM_LOW)
        `uvm_info(get_type_name(), $sformatf("  Data integrity priority mode: %s", data_integrity_priority ? "ENABLED" : "DISABLED"), UVM_LOW)
        `uvm_info(get_type_name(), $sformatf("  Level mismatch tolerance: %s", level_mismatch_tolerance ? "ENABLED" : "DISABLED"), UVM_LOW)
        `uvm_info(get_type_name(), $sformatf("  Underflow tolerance: %s", underflow_tolerance ? "ENABLED" : "DISABLED"), UVM_LOW)
        `uvm_info(get_type_name(), $sformatf("  Underflow tolerance count: %d", underflow_tolerance_count), UVM_LOW)
        `uvm_info(get_type_name(), $sformatf("  Write count tolerance: %s", write_count_tolerance ? "ENABLED" : "DISABLED"), UVM_LOW)
        `uvm_info(get_type_name(), $sformatf("  Write count tolerance count: %d", write_count_tolerance_count), UVM_LOW)
        `uvm_info(get_type_name(), $sformatf("  Reset scenario mode: %s", reset_scenario_active ? "ENABLED" : "DISABLED"), UVM_LOW)
        `uvm_info(get_type_name(), $sformatf("  Reset tolerance count: %d", reset_tolerance_count), UVM_LOW)
        if (error_count == 0) begin
            `uvm_info(get_type_name(), "Scoreboard: All checks passed!", UVM_LOW)
        end else begin
            `uvm_error(get_type_name(), $sformatf("Scoreboard: %d errors detected", error_count))
        end
    endfunction
    
    // Function to control data integrity priority settings
    function void set_data_integrity_priority(bit enable);
        data_integrity_priority = enable;
        `uvm_info(get_type_name(), $sformatf("Data integrity priority mode: %s", enable ? "ENABLED" : "DISABLED"), UVM_MEDIUM)
    endfunction
    
    // Function to control level mismatch tolerance
    function void set_level_mismatch_tolerance(bit enable);
        level_mismatch_tolerance = enable;
        `uvm_info(get_type_name(), $sformatf("Level mismatch tolerance: %s", enable ? "ENABLED" : "DISABLED"), UVM_MEDIUM)
    endfunction
    
    // Function to control use of actual RTL state for prev tracking
    function void set_use_actual_rtl_state(bit enable);
        use_actual_rtl_state = enable;
        `uvm_info(get_type_name(), $sformatf("Use actual RTL state for prev tracking: %s", enable ? "ENABLED" : "DISABLED"), UVM_MEDIUM)
    endfunction
    
    // Function to control underflow tolerance
    function void set_underflow_tolerance(bit enable);
        underflow_tolerance = enable;
        `uvm_info(get_type_name(), $sformatf("Underflow tolerance: %s", enable ? "ENABLED" : "DISABLED"), UVM_MEDIUM)
    endfunction
    
    // Function to control write count tolerance
    function void set_write_count_tolerance(bit enable);
        write_count_tolerance = enable;
        `uvm_info(get_type_name(), $sformatf("Write count tolerance: %s", enable ? "ENABLED" : "DISABLED"), UVM_MEDIUM)
    endfunction
    
    // Function to set reset scenario mode
    function void set_reset_scenario_mode(bit enable);
        reset_scenario_active = enable;
        `uvm_info(get_type_name(), $sformatf("Reset scenario mode: %s", enable ? "ENABLED" : "DISABLED"), UVM_MEDIUM)
    endfunction
    
    // Function to get data integrity statistics
    function void get_data_integrity_stats(output int total_ops, output int sim_ops, output int errors);
        total_ops = write_count + read_count;
        sim_ops = simultaneous_operation_count;
        errors = error_count;
    endfunction
    
    // Function to configure SOFT_RESET parameter
    function void set_soft_reset_param(int value);
        SOFT_RESET_PARAM = value;
        `uvm_info(get_type_name(), $sformatf("SOFT_RESET parameter set to: %0d", SOFT_RESET_PARAM), UVM_MEDIUM)
    endfunction
    
    // Function to configure SYNC_STAGE parameter
    function void set_sync_stage_param(int value);
        SYNC_STAGE_PARAM = value;
        `uvm_info(get_type_name(), $sformatf("SYNC_STAGE parameter set to: %0d", SYNC_STAGE_PARAM), UVM_MEDIUM)
    endfunction
    
    // Function to get current parameter values
    function void get_parameters(output int soft_reset, output int sync_stage);
        soft_reset = SOFT_RESET_PARAM;
        sync_stage = SYNC_STAGE_PARAM;
    endfunction
    
    // Function to calculate synchronization delay based on SYNC_STAGE
    function int get_sync_delay();
        // SYNC_STAGE determines the number of flip-flops in the synchronizer
        // For SYNC_STAGE=2: 2 flip-flops = 2 clock cycles delay
        // For SYNC_STAGE=3: 3 flip-flops = 3 clock cycles delay
        return SYNC_STAGE_PARAM;
    endfunction
    
    // Function to determine soft reset behavior based on SOFT_RESET parameter
    function void determine_soft_reset_behavior(output bit write_reset, output bit read_reset);
        case (SOFT_RESET_PARAM)
            0: begin
                // SOFT_RESET=0: No soft reset functionality
                write_reset = 0;
                read_reset = 0;
            end
            1: begin
                // SOFT_RESET=1: Read domain reset only
                write_reset = 0;
                read_reset = 1;
            end
            2: begin
                // SOFT_RESET=2: Write domain reset only
                write_reset = 1;
                read_reset = 0;
            end
            3: begin
                // SOFT_RESET=3: Both domains reset
                write_reset = 1;
                read_reset = 1;
            end
            default: begin
                // Default to no reset
                write_reset = 0;
                read_reset = 0;
            end
        endcase
    endfunction
    
    // Function to get human-readable soft reset description
    function string get_soft_reset_description();
        case (SOFT_RESET_PARAM)
            0: return "No soft reset functionality";
            1: return "Read domain reset only";
            2: return "Write domain reset only";
            3: return "Both domains reset";
            default: return "Unknown";
        endcase
    endfunction
endclass